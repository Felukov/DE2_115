library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity pit_counter is
    port (
        clk             : in std_logic;
        resetn          : in std_logic

    );
end entity pit_counter;

architecture rtl of pit_counter is

begin



end architecture;