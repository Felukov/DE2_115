
-- Copyright (C) 2022, Konstantin Felukov
-- All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- * Redistributions of source code must retain the above copyright notice, this
--   list of conditions and the following disclaimer.
--
-- * Redistributions in binary form must reproduce the above copyright notice,
--   this list of conditions and the following disclaimer in the documentation
--   and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
-- SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
-- CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
-- OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
-- OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.cpu86_types.all;

entity cpu86_bpu is
    port (
        clk                         : in std_logic;
        resetn                      : in std_logic;

        s_axis_instr_tvalid         : in std_logic;
        s_axis_instr_tready         : out std_logic;
        s_axis_instr_tdata          : in decoded_instr_t;
        s_axis_instr_tuser          : in user_t;

        m_axis_instr_tvalid         : out std_logic;
        m_axis_instr_tready         : in std_logic;
        m_axis_instr_tdata          : out decoded_instr_t;
        m_axis_instr_tuser          : out user_t;

        s_axis_jump_tvalid          : in std_logic;
        s_axis_jump_tdata           : in cpu86_jump_t;

        m_axis_jump_tvalid          : out std_logic;
        m_axis_jump_tdata           : out std_logic_vector(31 downto 0)
    );
end entity cpu86_bpu;

architecture rtl of cpu86_bpu is

    constant BPU_ITEM_CNT           : natural := 8;

    type bpu_item_t is record
        valid                       : std_logic;
        saturated_cnt               : natural range 0 to 3;
        inst_cs                     : std_logic_vector(15 downto 0);
        inst_ip                     : std_logic_vector(15 downto 0);
        jump_cs                     : std_logic_vector(15 downto 0);
        jump_ip                     : std_logic_vector(15 downto 0);
    end record;

    type bpu_items_t is array (natural range 0 to BPU_ITEM_CNT-1) of bpu_item_t;

    signal instr_s_tvalid           : std_logic;
    signal instr_s_tready           : std_logic;
    signal instr_s_tdata            : decoded_instr_t;
    signal instr_s_tuser            : user_t;

    signal instr_m_tvalid           : std_logic;
    signal instr_m_tready           : std_logic;
    signal instr_m_tdata            : decoded_instr_t;
    signal instr_m_tuser            : user_t;

    signal jump_s_tvalid            : std_logic;
    signal jump_s_tdata             : cpu86_jump_t;
    signal jump_m_tvalid            : std_logic;
    signal jump_m_tdata             : std_logic_vector(31 downto 0);

    signal bpu_items                : bpu_items_t;
    signal bpu_wr_valid             : std_logic;
    signal bpu_wr_idx               : natural range 0 to BPU_ITEM_CNT-1;
    signal bpu_rd_idx               : natural range 0 to BPU_ITEM_CNT-1;
    signal bpu_item_wr_hit          : std_logic_vector(BPU_ITEM_CNT-1 downto 0);
    signal bpu_item_wr_hit_any      : std_logic;

    signal bpu_item_rd_hit          : std_logic_vector(BPU_ITEM_CNT-1 downto 0);
    signal bpu_item_rd_hit_any      : std_logic;
    signal bpu_item_rd_hit_idx      : natural range 0 to BPU_ITEM_CNT-1;

    signal next_free_bpu_item_idx   : natural range 0 to BPU_ITEM_CNT-1;

    signal jump_pass                : std_logic;

begin
    -- i/o assigns
    instr_s_tvalid      <= s_axis_instr_tvalid;
    s_axis_instr_tready <= instr_s_tready;
    instr_s_tdata       <= s_axis_instr_tdata;
    instr_s_tuser       <= s_axis_instr_tuser;

    m_axis_instr_tvalid <= instr_m_tvalid;
    instr_m_tready      <= m_axis_instr_tready;
    m_axis_instr_tdata  <= instr_m_tdata;
    m_axis_instr_tuser  <= instr_m_tuser;

    jump_s_tvalid       <= s_axis_jump_tvalid;
    jump_s_tdata        <= s_axis_jump_tdata;

    m_axis_jump_tvalid  <= jump_m_tvalid;
    m_axis_jump_tdata   <= jump_m_tdata;

    -- assigns
    instr_s_tready      <= '1' when jump_s_tvalid = '0' and jump_m_tvalid = '0' and (instr_m_tvalid = '0' or (instr_m_tvalid = '1' and instr_m_tready = '1')) else '0';

    jump_pass           <= '1' when instr_s_tdata.op = BRANCH or instr_s_tdata.op = RET else '0';

    -- forwarding instruction
    process (clk) begin
        if rising_edge(clk) then
            -- resettable logic
            if resetn = '0' then
                instr_m_tvalid <= '0';
            else
                if (jump_s_tvalid = '1' and jump_s_tdata.mismatch = '1') then
                    instr_m_tvalid <= '0';
                elsif (instr_s_tvalid = '1' and instr_s_tready = '1') then
                    instr_m_tvalid <= '1';
                elsif (instr_m_tready = '1') then
                    instr_m_tvalid <= '0';
                end if;
            end if;

            --without reset
            if (instr_s_tvalid = '1' and instr_s_tready = '1') then
                if (bpu_item_rd_hit_any = '1' and
                    bpu_items(bpu_item_rd_hit_idx).saturated_cnt > 1 and
                    jump_pass = '1') then
                    instr_m_tdata.bpu_taken <= '1';
                else
                    instr_m_tdata.bpu_taken <= '0';
                end if;

                if (bpu_item_rd_hit_any = '1') then
                    instr_m_tdata.bpu_first <= '0';
                else
                    instr_m_tdata.bpu_first <= '1';
                end if;

                instr_m_tdata.bpu_taken_cs  <= bpu_items(bpu_item_rd_hit_idx).jump_cs;
                instr_m_tdata.bpu_taken_ip  <= bpu_items(bpu_item_rd_hit_idx).jump_ip;

                instr_m_tdata.op            <= instr_s_tdata.op;
                instr_m_tdata.code          <= instr_s_tdata.code;
                instr_m_tdata.w             <= instr_s_tdata.w;
                instr_m_tdata.dir           <= instr_s_tdata.dir;
                instr_m_tdata.ea            <= instr_s_tdata.ea;
                instr_m_tdata.dreg          <= instr_s_tdata.dreg;
                instr_m_tdata.dmask         <= instr_s_tdata.dmask;
                instr_m_tdata.sreg          <= instr_s_tdata.sreg;
                instr_m_tdata.smask         <= instr_s_tdata.smask;
                instr_m_tdata.data          <= instr_s_tdata.data;
                instr_m_tdata.disp          <= instr_s_tdata.disp;
                instr_m_tdata.fl            <= instr_s_tdata.fl;
                instr_m_tdata.imm8          <= instr_s_tdata.imm8;
                instr_m_tdata.wait_ax       <= instr_s_tdata.wait_ax;
                instr_m_tdata.wait_bx       <= instr_s_tdata.wait_bx;
                instr_m_tdata.wait_cx       <= instr_s_tdata.wait_cx;
                instr_m_tdata.wait_dx       <= instr_s_tdata.wait_dx;
                instr_m_tdata.wait_bp       <= instr_s_tdata.wait_bp;
                instr_m_tdata.wait_si       <= instr_s_tdata.wait_si;
                instr_m_tdata.wait_di       <= instr_s_tdata.wait_di;
                instr_m_tdata.wait_sp       <= instr_s_tdata.wait_sp;
                instr_m_tdata.wait_ds       <= instr_s_tdata.wait_ds;
                instr_m_tdata.wait_es       <= instr_s_tdata.wait_es;
                instr_m_tdata.wait_ss       <= instr_s_tdata.wait_ss;
                instr_m_tdata.wait_fl       <= instr_s_tdata.wait_fl;
                instr_m_tdata.lock_fl       <= instr_s_tdata.lock_fl;
                instr_m_tdata.lock_sreg     <= instr_s_tdata.lock_sreg;
                instr_m_tdata.lock_dreg     <= instr_s_tdata.lock_dreg;
                instr_m_tdata.lock_ax       <= instr_s_tdata.lock_ax;
                instr_m_tdata.lock_sp       <= instr_s_tdata.lock_sp;
                instr_m_tdata.lock_si       <= instr_s_tdata.lock_si;
                instr_m_tdata.lock_di       <= instr_s_tdata.lock_di;
                instr_m_tdata.lock_ds       <= instr_s_tdata.lock_ds;
                instr_m_tdata.lock_es       <= instr_s_tdata.lock_es;
                instr_m_tdata.lock_all      <= instr_s_tdata.lock_all;

                instr_m_tuser               <= instr_s_tuser;
            end if;
        end if;
    end process;

    -- driving jump
    jump_proc: process (clk) begin
        if rising_edge(clk) then
            -- resettable logic
            if resetn = '0' then
                jump_m_tvalid <= '0';
            else
                if ((jump_s_tvalid = '1' and jump_s_tdata.mismatch = '1') or
                    (instr_s_tvalid = '1' and instr_s_tready = '1' and instr_s_tdata.op = JMPU  and instr_s_tdata.code(3) = '0') or
                    (instr_s_tvalid = '1' and instr_s_tready = '1' and instr_s_tdata.op = JCALL and instr_s_tdata.code(3) = '0') or
                    (instr_s_tvalid = '1' and instr_s_tready = '1' and bpu_item_rd_hit_any = '1' and bpu_items(bpu_item_rd_hit_idx).saturated_cnt > 1 and jump_pass = '1'))
                then
                    jump_m_tvalid <= '1';
                else
                    jump_m_tvalid <= '0';
                end if;
            end if;

            -- without reset
            if (jump_s_tvalid = '1' and jump_s_tdata.mismatch = '1') then
                jump_m_tdata(31 downto 16) <= jump_s_tdata.jump_cs;
                jump_m_tdata(15 downto 0)  <= jump_s_tdata.jump_ip;
            elsif (instr_s_tvalid = '1' and instr_s_tready = '1' and (instr_s_tdata.op = JMPU or instr_s_tdata.op = JCALL)) then
                if (instr_s_tdata.code = JMP_PTR16_16 or instr_s_tdata.code = CALL_PTR16_16) then
                    jump_m_tdata(31 downto 16) <= instr_s_tdata.data;
                    jump_m_tdata(15 downto 0)  <= instr_s_tdata.disp;
                else
                    jump_m_tdata(31 downto 16) <= instr_s_tuser(31 downto 16);
                    jump_m_tdata(15 downto 0)  <= std_logic_vector(unsigned(instr_s_tuser(15 downto 0)) + unsigned(instr_s_tdata.disp));
                end if;
            elsif (instr_s_tvalid = '1' and instr_s_tready = '1') then
                jump_m_tdata(31 downto 16) <= bpu_items(bpu_item_rd_hit_idx).jump_cs;
                jump_m_tdata(15 downto 0)  <= bpu_items(bpu_item_rd_hit_idx).jump_ip;
            end if;
        end if;
    end process;

    bpu_item_wr_hit_gen : for i in 0 to BPU_ITEM_CNT-1 generate

        bpu_item_wr_hit(i) <= '1' when (bpu_items(i).valid = '1' and
            bpu_items(i).inst_cs = jump_s_tdata.inst_cs and
            bpu_items(i).inst_ip = jump_s_tdata.inst_ip)
        else '0';

    end generate;

    bpu_item_wr_hit_any <= '1' when bpu_item_wr_hit /= "00000000" else '0';

    process (all) begin
        for i in 0 to BPU_ITEM_CNT-1 loop

            if (bpu_items(i).valid = '1' and
                bpu_items(i).inst_cs = instr_s_tuser(USER_T_CS) and
                bpu_items(i).inst_ip = instr_s_tuser(USER_T_IP))
            then
                bpu_item_rd_hit(i) <= '1';
            else
                bpu_item_rd_hit(i) <= '0';
            end if;

        end loop;

        bpu_item_rd_hit_any <= '0';
        bpu_item_rd_hit_idx <= 0;
        for i in 0 to BPU_ITEM_CNT-1 loop
            if (bpu_item_rd_hit(i) = '1') then
                bpu_item_rd_hit_any <= '1';
                bpu_item_rd_hit_idx <= i;
            end if;
        end loop;

    end process;

    process (clk) begin
        if rising_edge(clk) then
            -- Resettable logic
            if resetn = '0' then
                for i in 0 to BPU_ITEM_CNT-1 loop
                    bpu_items(i).valid <= '0';
                end loop;
            else

                for i in 0 to BPU_ITEM_CNT-1 loop
                    if (jump_s_tvalid = '1' and jump_s_tdata.bypass = '0' and ((bpu_item_wr_hit(i) = '1') or (bpu_item_wr_hit_any = '0' and i = next_free_bpu_item_idx))) then
                        bpu_items(i).valid <= '1';
                    end if;
                end loop;

            end if;

            -- Without reset
            for i in 0 to BPU_ITEM_CNT-1 loop
                if (jump_s_tvalid = '1' and jump_s_tdata.bypass = '0' and ((bpu_item_wr_hit(i) = '1') or (bpu_item_wr_hit_any = '0' and i = next_free_bpu_item_idx))) then
                    bpu_items(i).inst_cs <= jump_s_tdata.inst_cs;
                    bpu_items(i).inst_ip <= jump_s_tdata.inst_ip;

                    if (jump_s_tdata.taken = '1') then
                        bpu_items(i).jump_cs <= jump_s_tdata.jump_cs;
                        bpu_items(i).jump_ip <= jump_s_tdata.jump_ip;
                    end if;

                    if (jump_s_tdata.first = '1') then
                        if (jump_s_tdata.taken = '1') then
                            bpu_items(i).saturated_cnt <= 1;
                        else
                            bpu_items(i).saturated_cnt <= 0;
                        end if;
                    else
                        if (jump_s_tdata.taken = '1' and bpu_items(i).saturated_cnt < 3) then
                            bpu_items(i).saturated_cnt <= bpu_items(i).saturated_cnt + 1;
                        elsif (jump_s_tdata.taken = '0' and bpu_items(i).saturated_cnt > 0) then
                            bpu_items(i).saturated_cnt <= bpu_items(i).saturated_cnt - 1;
                        end if;
                    end if;

                end if;
            end loop;

        end if;

    end process;

    process (clk) begin
        if rising_edge(clk) then
            if resetn = '0' then
                next_free_bpu_item_idx <= 0;
            else
                if (jump_s_tvalid = '1' and jump_s_tdata.bypass = '0' and bpu_item_wr_hit_any = '0') then
                    next_free_bpu_item_idx <= (next_free_bpu_item_idx + 1) mod BPU_ITEM_CNT;
                end if;
            end if;
        end if;
    end process;

end architecture;
